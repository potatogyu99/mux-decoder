module decoder_3to8 (
    input wire [2:0] in,  // 3비트 입력
    output reg [7:0] out  // 8개의 출력
);

always @(*)
begin
    case(in)
        3'b000: out = 8'b10000000; // 입력이 000이면 첫 번째 출력이 활성화됩니다.
        3'b001: out = 8'b01000000; // 입력이 001이면 두 번째 출력이 활성화됩니다.
        3'b010: out = 8'b00100000; // 입력이 010이면 세 번째 출력이 활성화됩니다.
        3'b011: out = 8'b00010000; // 입력이 011이면 네 번째 출력이 활성화됩니다.
        3'b100: out = 8'b00001000; // 입력이 100이면 다섯 번째 출력이 활성화됩니다.
        3'b101: out = 8'b00000100; // 입력이 101이면 여섯 번째 출력이 활성화됩니다.
        3'b110: out = 8'b00000010; // 입력이 110이면 일곱 번째 출력이 활성화됩니다.
        3'b111: out = 8'b00000001; // 입력이 111이면 여덟 번째 출력이 활성화됩니다.
        default: out = 8'b00000000; // 그 외의 경우 모든 출력이 비활성화됩니다.
    endcase
end

endmodule
